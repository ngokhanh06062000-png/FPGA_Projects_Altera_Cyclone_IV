module inv 
(
input logic [3:0] a,	// a[3:0] - 4-битная шина, биты от старшего к младшему так: a[3] a[2] a[1] a[0]
						// Это - little endian (младший бит имеет наименьший битовый номер)
						// Если a[0:3] тогда порядок битов от старшего к младшему как: a[0] a[1] a[2] a[3] 
						// Это - big endian
output logic [3:0] y
);

	assign y = ~a;

endmodule