module testbench1();
	logic a, b, c, y;
	
	// задание (определение) тестируемого устройства
	sillyfunction dut(a, b, c, y);
	
	// активировать входы пошагово с интервалом
	initial begin
		a = 0; b = 0; c = 0; 	#10;
		c = 1; 					#10;
		b = 1; c = 0;			#10;
		c = 1;					#10;
		a = 1; b = 0; c = 0;	#10;
		c = 1;					#10;
		b = 1; c = 0;			#10;
		c = 1;					#10;
	end
endmodule
/*
Оператор 'initial' выполняет содержащиеся в нем операторы в нулевой момент времени моделирования
в данном случае он подает на входы набор 000, 
ждет 10 единиц времени. Затем 001 и ждет ещё 10 единиц времени...

Оператор 'initial' должен быть использовать в тестбенчах для моделирования
а не в модулях, из которых будет синтезирована аппаратура
*/