/* Регистр */
module flop 
(
input logic 		clk,
input logic [3:0]	  d,
output logic [3:0]    q
);

	always_ff @(posedge clk)
		q <= d; 		// q принимает значение d
/*
		<= - неблокирующее присваивание, 
		используемый внутри оператора 'always' вместо 'assign'
		Так как операторы 'always' можно использовать для создания триггеров, защелок или комбинационной логики
 		Для избежания нежелательных ошибок, введены в Systemverilog:
		1) always_ff - синтез триггеров и позволять выдавать предупреждение
		инструментальной среде в противном случае
		2) always_latch - 
		3) always_comb - 
*/
endmodule