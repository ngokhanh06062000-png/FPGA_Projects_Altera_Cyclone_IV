module tristate 
(
input logic [3:0] a,
input logic 	  en,
output tri  [3:0] y  		// tri - тристабильная шина
);
/* 
logic - имеет только один драйвер
tri - может иметь несколько драйвер (Есть 2 применяемых типа tri и tri-reg)
Обычно один драйвер в сети активен в конкретный момент времени, 
если ни один из драйверов не активирован то tri = z - высокоимпедансное состояние 
и tri-reg = предыдущее значение
*/
	assign y = en ? a : 4'bz;

/* Манипуляция с битами */
/*
	assign y = {c[2:1], {3{d[0]}}, c[0], 3'b101};
	
	// y = c[2]c[1]d[0]d[0]d[0]c[0]101 
*/

endmodule

