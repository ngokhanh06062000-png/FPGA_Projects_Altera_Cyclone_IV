module inv
(
input logic [3:0]  a,
output logic [3:0] y
);

	always_comb		// 'always_comb' реагирует выражение внутри always каждый раз
					//  когда изменяется любой из сигналов правой части '<=' или '='
		y = ~a;		//  блокирующее присваивание
	/*
	В операторе 'always'
	Знак '=' - блокирующее
	Знак '<=' - неблокирующее присваивание (или одновременное)
	
	Не путайте эти присваивания с непрерывным присваиванием 
	с помощью оператора 'assign'
	'assign' используется вне операторов 'always' и тоже одновременное вычисляются 
	*/

endmodule